module frewsave(input A0,input CS1,
				input [15:0] Data_In
					);